library verilog;
use verilog.vl_types.all;
entity maior_vlg_vec_tst is
end maior_vlg_vec_tst;
