library verilog;
use verilog.vl_types.all;
entity subtracao_vlg_vec_tst is
end subtracao_vlg_vec_tst;
